`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//------------------------------------------------------------------------------------
//------------------------------------------------------------------------------------
//------------------------------------------------------------------------------------
// Create Date: 02/25/2020 11:40:30 AM
// Module Name: RCANew
// Project Name: Milestone #2
// Author:  Yasmin Elwazir  900161056
//          Donia Ghazy     900172124
//          Yousef Elwazir  900161060
// Description: Ripple Carry Adder with N=32 bits
// Change History:
//                  Last modified 19/04/2020
//------------------------------------------------------------------------------------
//------------------------------------------------------------------------------------
//------------------------------------------------------------------------------------



module RCANew #(parameter N=32) (input [N-1:0] A, input [N-1:0] B, output [N-1:0] C );


wire [N:0] carries;
assign carries[0]=0;

genvar i;
generate
for( i=0 ; i<32;i=i+1)
FullAdderNew adder( A[i],B[i],carries[i],C[i],carries[i+1]);
endgenerate



endmodule


