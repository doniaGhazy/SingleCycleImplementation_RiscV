`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//------------------------------------------------------------------------------------
//------------------------------------------------------------------------------------
//------------------------------------------------------------------------------------
// Create Date: 02/18/2020 11:29:50 AM
// Module Name: DFlipFlop
// Project Name: Milestone #2
// Author:  Yasmin Elwazir  900161056
//          Donia Ghazy     900172124
//          Yousef Elwazir  900161060
// Description: DFlipFlop
// Change History:
//                  Last Modified 19/04/2020
//------------------------------------------------------------------------------------
//------------------------------------------------------------------------------------
//------------------------------------------------------------------------------------


module DFlipFlop      (input clk, input rst, input D, output reg Q); 
 
    always @ (posedge clk or posedge rst)  
   if (!rst) begin    
     Q <= 1'b0;   
  end  else begin    
     Q <= D;   
  end 
endmodule 


